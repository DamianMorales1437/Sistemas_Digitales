//Compuerta XOR

module Compuerta_xor(
	input A,
	input B,
	output F
	);

assign F = A ^ B;
endmodule
