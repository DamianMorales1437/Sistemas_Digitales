module primera_funcion(
//entradas y salidas
//modo tipo ancho nombre
 input A,B,
 output F
);
assign F=~A|B;
endmodule