module comparador(
    input [2:0] A, B,
	output F    
);
// DECLARACIÓN DE VARIABLES

// ==========================
// DESCRIPCIÓN DEL CIRCUITO
assign F = A > B;

endmodule 