//Compuerta AND

module Compuerta_and(
	input A,
	input B,
	output F
	);

assign F = A & B;
endmodule
