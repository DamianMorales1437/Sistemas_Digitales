module sum(
   input [2:0] A,B,
   output [3:0] F    
);
// DECLARACIÓN DE VARIABLES

// ==========================
// DESCRIPCIÓN DEL CIRCUITO
assign F = A + B;

endmodule 