`timescale 1ns / 1ps
//Codificador
module deco(
input [3:0] S,
input [8:0] C50,C20,C10,C5,
output reg [8:0] F
);

always @(*)
        case (S)
            4'b1000 : begin
	            case({C50})	            
	            9'd0: F = 9'b000000000;
	            9'd1: F = 9'b000000001;
	            9'd2: F = 9'b000000011;
	            9'd3: F = 9'b000000111;
	            9'd4: F = 9'b000001111;
	            9'd5: F = 9'b000011111;
	            9'd6: F = 9'b000111111;
	            9'd7: F = 9'b001111111;
	            9'd8: F = 9'b011111111;	
	            endcase
                      end
            4'b0100: begin
	            case({C20})	            
	            9'd0: F = 9'b000000000;
	            9'd1: F = 9'b000000001;
	            9'd2: F = 9'b000000011;
	            9'd3: F = 9'b000000111;
	            9'd4: F = 9'b000001111;
	            9'd5: F = 9'b000011111;
	            9'd6: F = 9'b000111111;
	            9'd7: F = 9'b001111111;
	            9'd8: F = 9'b011111111;	            
	            endcase
                      end
             4'b0010: begin
                case({C10})                
	            9'd0: F = 9'b000000000;
	            9'd1: F = 9'b000000001;
	            9'd2: F = 9'b000000011;
	            9'd3: F = 9'b000000111;
	            9'd4: F = 9'b000001111;
	            9'd5: F = 9'b000011111;
	            9'd6: F = 9'b000111111;
	            9'd7: F = 9'b001111111;
	            9'd8: F = 9'b011111111;	
                endcase
                      end
			 4'b0001: begin
                case({C5})                
	            9'd0: F = 9'b000000000;
	            9'd1: F = 9'b000000001;
	            9'd2: F = 9'b000000011;
	            9'd3: F = 9'b000000111;
	            9'd4: F = 9'b000001111;
	            9'd5: F = 9'b000011111;
	            9'd6: F = 9'b000111111;
	            9'd7: F = 9'b001111111;
	            9'd8: F = 9'b011111111;	
                endcase     
                      end
	    endcase 				  
endmodule
