module NombreModulo_Labsland
(   // Utilizar los nombres de los puertos 
    // indicados en la documentación en LabsLand
    // INPUT: SW - KEY - CLOCK_50
    // OUTPUT: LEDR - HEXn
    
);
// ===============================================
// CONEXIÓN DEL CIRCUITO QUE SE QUIERE IMPLEMENTAR
NombreCircuito  etiqueta(
  .entrada_circuito(puerto_labsland),
  .entrada_circuito(puerto_labsland),
  .salida_circuito(puerto_labsland)
  .salida_circuito(puerto_labsland)
);
// -----------------------------------------------
endmodule