//Compuerta NOT

module Compuerta_not(
	input A,
	output F
	);

assign F = ~A;
endmodule
