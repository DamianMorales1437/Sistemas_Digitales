module NombreModuloCircuito
(   // ENTRADAS y SALIDAS
    
    
);
// = = = = = = = = = = = = =
// DECLARACIÓN DE VARIABLES


// -------------------------


// = = = = = = = = = = = = =
// DESCRIPCIÓN DEL CIRCUITO


// -------------------------
endmodule 