//Compuerta OR

module Compuerta_or(
	input A,
	input B,
	output F
	);

assign F = A | B;
endmodule
